/*Program for driving a seven segment display
January 18,2021
Code by G V V Sharma
Released under GNU GPL
*/

//declaring the blink module
module helloworldfpga(
                 output a,
                 output b,
                 output c,
             output d,
               output e,
              output f,
               output g

);

assign     a=1;
assign     b=0;
assign     c=0;
assign     d=1;
assign     e=1;
assign     f=1;
assign     g=1;
endmodule
//end of the module







